{"Level": "1", "Exp": "0", "Money": "0", "Target": "\u041e\u0442\u043c\u0435\u043d\u0438\u0442\u044c \u0434/\u0437"}